module Mult_Combinational(
    input [3:0] ABus, BBus,
    input [3:0] Areg, Breg, Preg,
    input [5:0] ps,
    input _192_, start,

    output _193_, _024_, 
    output [3:0] _000_, _001_, _002_,
    output ready,
    output [7:0] resultBus
);

  wire _003_;
  wire _004_;
  wire _005_;
  wire _006_;
  wire _007_;
  wire _008_;
  wire _009_;
  wire _010_;
  wire _011_;
  wire _012_;
  wire _013_;
  wire _014_;
  wire _015_;
  wire _016_;
  wire _017_;
  wire _018_;
  wire _019_;
  wire _020_;
  wire _021_;
  wire _022_;
  wire _023_;
  wire _025_;
  wire _026_;
  wire _027_;
  wire _028_;
  wire _029_;
  wire _030_;
  wire _031_;
  wire _032_;
  wire _033_;
  wire _034_;
  wire _035_;
  wire _036_;
  wire _037_;
  wire _038_;
  wire _039_;
  wire _040_;
  wire _041_;
  wire _042_;
  wire _043_;
  wire _044_;
  wire _045_;
  wire _046_;
  wire _047_;
  wire _048_;
  wire _049_;
  wire _050_;
  wire _051_;
  wire _052_;
  wire _053_;
  wire _054_;
  wire _055_;
  wire _056_;
  wire _057_;
  wire _058_;
  wire _059_;
  wire _060_;
  wire _061_;
  wire _062_;
  wire _063_;
  wire _064_;
  wire _065_;
  wire _066_;
  wire _067_;
  wire _068_;
  wire _069_;
  wire _070_;
  wire _071_;
  wire _072_;
  wire _073_;
  wire _074_;
  wire _075_;
  wire _076_;
  wire _077_;
  wire _078_;
  wire _079_;
  wire _080_;
  wire _081_;
  wire _082_;
  wire _083_;
  wire _084_;
  wire _085_;
  wire _086_;
  wire _087_;
  wire _088_;
  wire _089_;
  wire _090_;
  wire _091_;
  wire _092_;
  wire _093_;
  wire _094_;
  wire _095_;
  wire _096_;
  wire _097_;
  wire _098_;
  wire _099_;
  wire _100_;
  wire _101_;
  wire _102_;
  wire _103_;
  wire _104_;
  wire _105_;
  wire _106_;
  wire _107_;
  wire _108_;
  wire _109_;
  wire _110_;
  wire _111_;
  wire _112_;
  wire _113_;
  wire _114_;
  wire _115_;
  wire _116_;
  wire _117_;
  wire _118_;
  wire _119_;
  wire _120_;
  wire _121_;
  wire _122_;
  wire _123_;
  wire _124_;
  wire _125_;
  wire _126_;
  wire _127_;
  wire _128_;
  wire _129_;
  wire _130_;
  wire _131_;
  wire _132_;
  wire _133_;
  wire _134_;
  wire _135_;
  wire _136_;
  wire _137_;
  wire _138_;
  wire _139_;
  wire _140_;
  wire _141_;
  wire _142_;
  wire _143_;
  wire _144_;
  wire _145_;
  wire _146_;
  wire _147_;
  wire _148_;
  wire _149_;
  wire _150_;
  wire _151_;
  wire _152_;
  wire _153_;
  wire _154_;
  wire _155_;
  wire _156_;
  wire _157_;
  wire _158_;
  wire _159_;
  wire _160_;
  wire _161_;
  wire _162_;
  wire _163_;
  wire _164_;
  wire _165_;
  wire _166_;
  wire _167_;
  wire _168_;
  wire _169_;
  wire _170_;
  wire _171_;
  wire _172_;
  wire _173_;
  wire _174_;
  wire _175_;
  wire _176_;
  wire _177_;
  wire _178_;
  wire _179_;
  wire _180_;
  wire _181_;
  wire _182_;
  wire _183_;
  wire _184_;
  wire _185_;
  wire _186_;
  wire _187_;
  wire _188_;
  wire _189_;
  wire _190_;
  wire _191_;
  wire A0;
  wire initP;
  wire loadA;
  wire loadB;
  
  assign A0 = Areg[0];
  assign initP = ps[3];
  assign loadA = ps[3];
  assign loadB = ps[3];
  assign resultBus = { Preg, Areg };
  assign _109_ = start;
  assign _129_ = Preg[0];
  assign _165_ = ps[4];
  assign _182_ = ps[5];
  assign _062_ = ps[1];
  assign _071_ = ps[2];
  assign _095_ = Breg[1];
  assign _101_ = Areg[0];
  assign _103_ = Preg[1];
  assign _104_ = Breg[0];
  assign _105_ = ps[3];
  assign _107_ = Preg[2];
  assign _108_ = Breg[2];
  assign _113_ = Breg[3];
  assign _114_ = Preg[3];
  assign _134_ = BBus[0];
  assign _138_ = BBus[1];
  assign _142_ = BBus[2];
  assign _146_ = BBus[3];
  assign _150_ = Areg[1];
  assign _153_ = ABus[0];
  assign _157_ = Areg[2];
  assign _160_ = ABus[1];
  assign _164_ = Areg[3];
  assign _167_ = ABus[2];
  assign _173_ = ABus[3];
  assign _179_ = _192_;

  NOT _194_ (
    .A(_165_),
    .Y(_110_)
  );
  OR _195_ (
    .A(_179_),
    .B(_109_),
    .Y(_112_)
  );
  AND _196_ (
    .A(_112_),
    .B(_110_),
    .Y(_051_)
  );
  NOT _197_ (
    .A(_179_),
    .Y(_102_)
  );
  NOT _198_ (
    .A(_182_),
    .Y(_115_)
  );
  NOT _199_ (
    .A(_062_),
    .Y(_116_)
  );
  AND _200_ (
    .A(_116_),
    .B(_115_),
    .Y(_117_)
  );
  NOT _201_ (
    .A(_071_),
    .Y(_118_)
  );
  AND _202_ (
    .A(_118_),
    .B(_110_),
    .Y(_119_)
  );
  AND _203_ (
    .A(_119_),
    .B(_117_),
    .Y(_120_)
  );
  OR _204_ (
    .A(_062_),
    .B(_182_),
    .Y(_122_)
  );
  OR _205_ (
    .A(_071_),
    .B(_165_),
    .Y(_123_)
  );
  OR _206_ (
    .A(_123_),
    .B(_122_),
    .Y(_124_)
  );
  AND _207_ (
    .A(_124_),
    .B(_101_),
    .Y(_125_)
  );
  AND _208_ (
    .A(_125_),
    .B(_104_),
    .Y(_126_)
  );
  AND _209_ (
    .A(_126_),
    .B(_129_),
    .Y(_127_)
  );
  NOT _210_ (
    .A(_127_),
    .Y(_128_)
  );
  NOT _211_ (
    .A(_103_),
    .Y(_130_)
  );
  NOT _212_ (
    .A(_095_),
    .Y(_131_)
  );
  NOT _213_ (
    .A(_101_),
    .Y(_133_)
  );
  OR _214_ (
    .A(_120_),
    .B(_133_),
    .Y(_135_)
  );
  OR _215_ (
    .A(_135_),
    .B(_131_),
    .Y(_137_)
  );
  AND _216_ (
    .A(_137_),
    .B(_130_),
    .Y(_139_)
  );
  AND _217_ (
    .A(_125_),
    .B(_095_),
    .Y(_141_)
  );
  AND _218_ (
    .A(_141_),
    .B(_103_),
    .Y(_143_)
  );
  OR _219_ (
    .A(_143_),
    .B(_139_),
    .Y(_145_)
  );
  OR _220_ (
    .A(_145_),
    .B(_128_),
    .Y(_147_)
  );
  OR _221_ (
    .A(_141_),
    .B(_103_),
    .Y(_149_)
  );
  OR _222_ (
    .A(_137_),
    .B(_130_),
    .Y(_151_)
  );
  AND _223_ (
    .A(_151_),
    .B(_149_),
    .Y(_152_)
  );
  OR _224_ (
    .A(_152_),
    .B(_127_),
    .Y(_154_)
  );
  AND _225_ (
    .A(_154_),
    .B(_147_),
    .Y(_156_)
  );
  OR _226_ (
    .A(_156_),
    .B(_120_),
    .Y(_158_)
  );
  NOT _227_ (
    .A(_105_),
    .Y(_159_)
  );
  OR _228_ (
    .A(_124_),
    .B(_129_),
    .Y(_161_)
  );
  AND _229_ (
    .A(_161_),
    .B(_159_),
    .Y(_163_)
  );
  AND _230_ (
    .A(_163_),
    .B(_158_),
    .Y(_106_)
  );
  AND _231_ (
    .A(_152_),
    .B(_127_),
    .Y(_166_)
  );
  OR _232_ (
    .A(_166_),
    .B(_143_),
    .Y(_168_)
  );
  AND _233_ (
    .A(_125_),
    .B(_108_),
    .Y(_170_)
  );
  AND _234_ (
    .A(_170_),
    .B(_107_),
    .Y(_171_)
  );
  NOT _235_ (
    .A(_171_),
    .Y(_172_)
  );
  OR _236_ (
    .A(_170_),
    .B(_107_),
    .Y(_174_)
  );
  AND _237_ (
    .A(_174_),
    .B(_172_),
    .Y(_176_)
  );
  OR _238_ (
    .A(_176_),
    .B(_168_),
    .Y(_178_)
  );
  AND _239_ (
    .A(_147_),
    .B(_151_),
    .Y(_180_)
  );
  NOT _240_ (
    .A(_176_),
    .Y(_181_)
  );
  OR _241_ (
    .A(_181_),
    .B(_180_),
    .Y(_183_)
  );
  AND _242_ (
    .A(_183_),
    .B(_178_),
    .Y(_184_)
  );
  OR _243_ (
    .A(_184_),
    .B(_120_),
    .Y(_185_)
  );
  OR _244_ (
    .A(_124_),
    .B(_103_),
    .Y(_186_)
  );
  AND _245_ (
    .A(_186_),
    .B(_159_),
    .Y(_187_)
  );
  AND _246_ (
    .A(_187_),
    .B(_185_),
    .Y(_111_)
  );
  AND _247_ (
    .A(_183_),
    .B(_172_),
    .Y(_188_)
  );
  AND _248_ (
    .A(_125_),
    .B(_113_),
    .Y(_189_)
  );
  OR _249_ (
    .A(_189_),
    .B(_114_),
    .Y(_190_)
  );
  AND _250_ (
    .A(_189_),
    .B(_114_),
    .Y(_191_)
  );
  NOT _251_ (
    .A(_191_),
    .Y(_052_)
  );
  AND _252_ (
    .A(_052_),
    .B(_190_),
    .Y(_053_)
  );
  NOT _253_ (
    .A(_053_),
    .Y(_054_)
  );
  OR _254_ (
    .A(_054_),
    .B(_188_),
    .Y(_055_)
  );
  AND _255_ (
    .A(_176_),
    .B(_168_),
    .Y(_056_)
  );
  OR _256_ (
    .A(_056_),
    .B(_171_),
    .Y(_057_)
  );
  OR _257_ (
    .A(_053_),
    .B(_057_),
    .Y(_058_)
  );
  AND _258_ (
    .A(_058_),
    .B(_055_),
    .Y(_059_)
  );
  OR _259_ (
    .A(_059_),
    .B(_120_),
    .Y(_060_)
  );
  OR _260_ (
    .A(_124_),
    .B(_107_),
    .Y(_061_)
  );
  AND _261_ (
    .A(_061_),
    .B(_159_),
    .Y(_063_)
  );
  AND _262_ (
    .A(_063_),
    .B(_060_),
    .Y(_121_)
  );
  AND _263_ (
    .A(_053_),
    .B(_057_),
    .Y(_064_)
  );
  OR _264_ (
    .A(_191_),
    .B(_120_),
    .Y(_065_)
  );
  OR _265_ (
    .A(_065_),
    .B(_064_),
    .Y(_066_)
  );
  OR _266_ (
    .A(_124_),
    .B(_114_),
    .Y(_067_)
  );
  AND _267_ (
    .A(_067_),
    .B(_159_),
    .Y(_068_)
  );
  AND _268_ (
    .A(_068_),
    .B(_066_),
    .Y(_132_)
  );
  OR _269_ (
    .A(_105_),
    .B(_104_),
    .Y(_069_)
  );
  OR _270_ (
    .A(_134_),
    .B(_159_),
    .Y(_070_)
  );
  AND _271_ (
    .A(_070_),
    .B(_069_),
    .Y(_136_)
  );
  OR _272_ (
    .A(_105_),
    .B(_095_),
    .Y(_072_)
  );
  OR _273_ (
    .A(_138_),
    .B(_159_),
    .Y(_073_)
  );
  AND _274_ (
    .A(_073_),
    .B(_072_),
    .Y(_140_)
  );
  OR _275_ (
    .A(_108_),
    .B(_105_),
    .Y(_074_)
  );
  OR _276_ (
    .A(_142_),
    .B(_159_),
    .Y(_075_)
  );
  AND _277_ (
    .A(_075_),
    .B(_074_),
    .Y(_144_)
  );
  OR _278_ (
    .A(_113_),
    .B(_105_),
    .Y(_076_)
  );
  OR _279_ (
    .A(_146_),
    .B(_159_),
    .Y(_077_)
  );
  AND _280_ (
    .A(_077_),
    .B(_076_),
    .Y(_148_)
  );
  AND _281_ (
    .A(_120_),
    .B(_101_),
    .Y(_078_)
  );
  AND _282_ (
    .A(_124_),
    .B(_150_),
    .Y(_079_)
  );
  OR _283_ (
    .A(_079_),
    .B(_078_),
    .Y(_080_)
  );
  AND _284_ (
    .A(_080_),
    .B(_159_),
    .Y(_081_)
  );
  AND _285_ (
    .A(_153_),
    .B(_105_),
    .Y(_082_)
  );
  OR _286_ (
    .A(_082_),
    .B(_081_),
    .Y(_155_)
  );
  AND _287_ (
    .A(_120_),
    .B(_150_),
    .Y(_083_)
  );
  AND _288_ (
    .A(_124_),
    .B(_157_),
    .Y(_084_)
  );
  OR _289_ (
    .A(_084_),
    .B(_083_),
    .Y(_085_)
  );
  AND _290_ (
    .A(_085_),
    .B(_159_),
    .Y(_086_)
  );
  AND _291_ (
    .A(_160_),
    .B(_105_),
    .Y(_087_)
  );
  OR _292_ (
    .A(_087_),
    .B(_086_),
    .Y(_162_)
  );
  AND _293_ (
    .A(_120_),
    .B(_157_),
    .Y(_088_)
  );
  AND _294_ (
    .A(_124_),
    .B(_164_),
    .Y(_089_)
  );
  OR _295_ (
    .A(_089_),
    .B(_088_),
    .Y(_090_)
  );
  AND _296_ (
    .A(_090_),
    .B(_159_),
    .Y(_091_)
  );
  AND _297_ (
    .A(_167_),
    .B(_105_),
    .Y(_092_)
  );
  OR _298_ (
    .A(_092_),
    .B(_091_),
    .Y(_169_)
  );
  OR _299_ (
    .A(_173_),
    .B(_159_),
    .Y(_093_)
  );
  OR _300_ (
    .A(_126_),
    .B(_129_),
    .Y(_094_)
  );
  AND _301_ (
    .A(_128_),
    .B(_124_),
    .Y(_096_)
  );
  AND _302_ (
    .A(_096_),
    .B(_094_),
    .Y(_097_)
  );
  AND _303_ (
    .A(_120_),
    .B(_164_),
    .Y(_098_)
  );
  OR _304_ (
    .A(_098_),
    .B(_105_),
    .Y(_099_)
  );
  OR _305_ (
    .A(_099_),
    .B(_097_),
    .Y(_100_)
  );
  AND _306_ (
    .A(_100_),
    .B(_093_),
    .Y(_175_)
  );
  AND _307_ (
    .A(_102_),
    .B(_109_),
    .Y(_177_)
  );


  assign _193_ = _051_;
  assign ready = ps[0];
  assign ps[0] = _102_;
  assign _002_[0] = _106_;
  assign _002_[1] = _111_;
  assign _002_[2] = _121_;
  assign _002_[3] = _132_;
  assign _001_[0] = _136_;
  assign _001_[1] = _140_;
  assign _001_[2] = _144_;
  assign _001_[3] = _148_;
  assign _000_[0] = _155_;
  assign _000_[1] = _162_;
  assign _000_[2] = _169_;
  assign _000_[3] = _175_;
  assign _024_ = _177_;

endmodule
