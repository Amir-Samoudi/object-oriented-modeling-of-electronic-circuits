module Mult_Combinational_Behavioral(
    input [3:0] ABus,
    input [3:0] BBus,
    input [3:0] Areg,
    input [3:0] Breg,
    input [3:0] Preg,
    input [5:0] ps,
    input _192_,
    input start,
    output _193_,
    output _024_, 
    output [3:0] _000_,
    output [3:0] _001_,
    output [3:0] _002_,
    output ready,
    output [7:0] resultBus
);
    assign _193_ = ((((_192_) | (start)) & (~((ps[4])))));
    assign _024_ = (((~((_192_))) & (start)));
    assign _000_[0] = ((((ABus[0]) & (ps[3])) | ((((((ps[2]) | (ps[4])) | ((ps[1]) | (ps[5]))) & (Areg[1])) | ((((~((ps[2]))) & (~((ps[4])))) & ((~((ps[1]))) & (~((ps[5]))))) & (Areg[0]))) & (~((ps[3]))))));
    assign _000_[1] = ((((ABus[1]) & (ps[3])) | ((((((ps[2]) | (ps[4])) | ((ps[1]) | (ps[5]))) & (Areg[2])) | ((((~((ps[2]))) & (~((ps[4])))) & ((~((ps[1]))) & (~((ps[5]))))) & (Areg[1]))) & (~((ps[3]))))));
    assign _000_[2] = ((((ABus[2]) & (ps[3])) | ((((((ps[2]) | (ps[4])) | ((ps[1]) | (ps[5]))) & (Areg[3])) | ((((~((ps[2]))) & (~((ps[4])))) & ((~((ps[1]))) & (~((ps[5]))))) & (Areg[2]))) & (~((ps[3]))))));
    assign _000_[3] = ((((((((~((ps[2]))) & (~((ps[4])))) & ((~((ps[1]))) & (~((ps[5]))))) & (Areg[3])) | (ps[3])) | (((~(((((((ps[2]) | (ps[4])) | ((ps[1]) | (ps[5]))) & (Areg[0])) & (Breg[0])) & (Preg[0])))) & (((ps[2]) | (ps[4])) | ((ps[1]) | (ps[5])))) & ((((((ps[2]) | (ps[4])) | ((ps[1]) | (ps[5]))) & (Areg[0])) & (Breg[0])) | (Preg[0])))) & ((ABus[3]) | (~((ps[3]))))));
    assign _001_[0] = ((((BBus[0]) | (~((ps[3])))) & ((ps[3]) | (Breg[0]))));
    assign _001_[1] = ((((BBus[1]) | (~((ps[3])))) & ((ps[3]) | (Breg[1]))));
    assign _001_[2] = ((((BBus[2]) | (~((ps[3])))) & ((Breg[2]) | (ps[3]))));
    assign _001_[3] = ((((BBus[3]) | (~((ps[3])))) & ((Breg[3]) | (ps[3]))));
    assign _002_[0] = (((((((ps[2]) | (ps[4])) | ((ps[1]) | (ps[5]))) | (Preg[0])) & (~((ps[3])))) & ((((((((((~((ps[2]))) & (~((ps[4])))) & ((~((ps[1]))) & (~((ps[5]))))) | (~((Areg[0])))) | (~((Breg[1])))) | (~((Preg[1])))) & ((((((ps[2]) | (ps[4])) | ((ps[1]) | (ps[5]))) & (Areg[0])) & (Breg[1])) | (Preg[1]))) | ((((((ps[2]) | (ps[4])) | ((ps[1]) | (ps[5]))) & (Areg[0])) & (Breg[0])) & (Preg[0]))) & ((((((((ps[2]) | (ps[4])) | ((ps[1]) | (ps[5]))) & (Areg[0])) & (Breg[1])) & (Preg[1])) | ((((((~((ps[2]))) & (~((ps[4])))) & ((~((ps[1]))) & (~((ps[5]))))) | (~((Areg[0])))) | (~((Breg[1])))) & (~((Preg[1]))))) | (~(((((((ps[2]) | (ps[4])) | ((ps[1]) | (ps[5]))) & (Areg[0])) & (Breg[0])) & (Preg[0])))))) | (((~((ps[2]))) & (~((ps[4])))) & ((~((ps[1]))) & (~((ps[5]))))))));
    assign _002_[1] = (((((((ps[2]) | (ps[4])) | ((ps[1]) | (ps[5]))) | (Preg[1])) & (~((ps[3])))) & ((((~((((((((ps[2]) | (ps[4])) | ((ps[1]) | (ps[5]))) & (Areg[0])) & (Breg[2])) | (Preg[2])) & (~(((((((ps[2]) | (ps[4])) | ((ps[1]) | (ps[5]))) & (Areg[0])) & (Breg[2])) & (Preg[2]))))))) | (((((((((ps[2]) | (ps[4])) | ((ps[1]) | (ps[5]))) & (Areg[0])) & (Breg[1])) & (Preg[1])) | ((((((~((ps[2]))) & (~((ps[4])))) & ((~((ps[1]))) & (~((ps[5]))))) | (~((Areg[0])))) | (~((Breg[1])))) & (~((Preg[1]))))) | (~(((((((ps[2]) | (ps[4])) | ((ps[1]) | (ps[5]))) & (Areg[0])) & (Breg[0])) & (Preg[0]))))) & ((((((~((ps[2]))) & (~((ps[4])))) & ((~((ps[1]))) & (~((ps[5]))))) | (~((Areg[0])))) | (~((Breg[1])))) | (~((Preg[1])))))) & ((((((((ps[2]) | (ps[4])) | ((ps[1]) | (ps[5]))) & (Areg[0])) & (Breg[2])) | (Preg[2])) & (~(((((((ps[2]) | (ps[4])) | ((ps[1]) | (ps[5]))) & (Areg[0])) & (Breg[2])) & (Preg[2]))))) | (((((((((~((ps[2]))) & (~((ps[4])))) & ((~((ps[1]))) & (~((ps[5]))))) | (~((Areg[0])))) | (~((Breg[1])))) | (~((Preg[1])))) & ((((((ps[2]) | (ps[4])) | ((ps[1]) | (ps[5]))) & (Areg[0])) & (Breg[1])) | (Preg[1]))) & ((((((ps[2]) | (ps[4])) | ((ps[1]) | (ps[5]))) & (Areg[0])) & (Breg[0])) & (Preg[0]))) | ((((((ps[2]) | (ps[4])) | ((ps[1]) | (ps[5]))) & (Areg[0])) & (Breg[1])) & (Preg[1]))))) | (((~((ps[2]))) & (~((ps[4])))) & ((~((ps[1]))) & (~((ps[5]))))))));
    assign _002_[2] = (((((((ps[2]) | (ps[4])) | ((ps[1]) | (ps[5]))) | (Preg[2])) & (~((ps[3])))) & (((((~(((((((ps[2]) | (ps[4])) | ((ps[1]) | (ps[5]))) & (Areg[0])) & (Breg[3])) & (Preg[3])))) & ((((((ps[2]) | (ps[4])) | ((ps[1]) | (ps[5]))) & (Areg[0])) & (Breg[3])) | (Preg[3]))) | (((((((((ps[2]) | (ps[4])) | ((ps[1]) | (ps[5]))) & (Areg[0])) & (Breg[2])) | (Preg[2])) & (~(((((((ps[2]) | (ps[4])) | ((ps[1]) | (ps[5]))) & (Areg[0])) & (Breg[2])) & (Preg[2]))))) & (((((((((~((ps[2]))) & (~((ps[4])))) & ((~((ps[1]))) & (~((ps[5]))))) | (~((Areg[0])))) | (~((Breg[1])))) | (~((Preg[1])))) & ((((((ps[2]) | (ps[4])) | ((ps[1]) | (ps[5]))) & (Areg[0])) & (Breg[1])) | (Preg[1]))) & ((((((ps[2]) | (ps[4])) | ((ps[1]) | (ps[5]))) & (Areg[0])) & (Breg[0])) & (Preg[0]))) | ((((((ps[2]) | (ps[4])) | ((ps[1]) | (ps[5]))) & (Areg[0])) & (Breg[1])) & (Preg[1])))) | ((((((ps[2]) | (ps[4])) | ((ps[1]) | (ps[5]))) & (Areg[0])) & (Breg[2])) & (Preg[2])))) & ((~(((~(((((((ps[2]) | (ps[4])) | ((ps[1]) | (ps[5]))) & (Areg[0])) & (Breg[3])) & (Preg[3])))) & ((((((ps[2]) | (ps[4])) | ((ps[1]) | (ps[5]))) & (Areg[0])) & (Breg[3])) | (Preg[3]))))) | (((~((((((((ps[2]) | (ps[4])) | ((ps[1]) | (ps[5]))) & (Areg[0])) & (Breg[2])) | (Preg[2])) & (~(((((((ps[2]) | (ps[4])) | ((ps[1]) | (ps[5]))) & (Areg[0])) & (Breg[2])) & (Preg[2]))))))) | (((((((((ps[2]) | (ps[4])) | ((ps[1]) | (ps[5]))) & (Areg[0])) & (Breg[1])) & (Preg[1])) | ((((((~((ps[2]))) & (~((ps[4])))) & ((~((ps[1]))) & (~((ps[5]))))) | (~((Areg[0])))) | (~((Breg[1])))) & (~((Preg[1]))))) | (~(((((((ps[2]) | (ps[4])) | ((ps[1]) | (ps[5]))) & (Areg[0])) & (Breg[0])) & (Preg[0]))))) & ((((((~((ps[2]))) & (~((ps[4])))) & ((~((ps[1]))) & (~((ps[5]))))) | (~((Areg[0])))) | (~((Breg[1])))) | (~((Preg[1])))))) & (~(((((((ps[2]) | (ps[4])) | ((ps[1]) | (ps[5]))) & (Areg[0])) & (Breg[2])) & (Preg[2]))))))) | (((~((ps[2]))) & (~((ps[4])))) & ((~((ps[1]))) & (~((ps[5]))))))));
    assign _002_[3] = (((((((ps[2]) | (ps[4])) | ((ps[1]) | (ps[5]))) | (Preg[3])) & (~((ps[3])))) & ((((((((ps[2]) | (ps[4])) | ((ps[1]) | (ps[5]))) & (Areg[0])) & (Breg[3])) & (Preg[3])) | (((~((ps[2]))) & (~((ps[4])))) & ((~((ps[1]))) & (~((ps[5])))))) | (((~(((((((ps[2]) | (ps[4])) | ((ps[1]) | (ps[5]))) & (Areg[0])) & (Breg[3])) & (Preg[3])))) & ((((((ps[2]) | (ps[4])) | ((ps[1]) | (ps[5]))) & (Areg[0])) & (Breg[3])) | (Preg[3]))) & (((((((((ps[2]) | (ps[4])) | ((ps[1]) | (ps[5]))) & (Areg[0])) & (Breg[2])) | (Preg[2])) & (~(((((((ps[2]) | (ps[4])) | ((ps[1]) | (ps[5]))) & (Areg[0])) & (Breg[2])) & (Preg[2]))))) & (((((((((~((ps[2]))) & (~((ps[4])))) & ((~((ps[1]))) & (~((ps[5]))))) | (~((Areg[0])))) | (~((Breg[1])))) | (~((Preg[1])))) & ((((((ps[2]) | (ps[4])) | ((ps[1]) | (ps[5]))) & (Areg[0])) & (Breg[1])) | (Preg[1]))) & ((((((ps[2]) | (ps[4])) | ((ps[1]) | (ps[5]))) & (Areg[0])) & (Breg[0])) & (Preg[0]))) | ((((((ps[2]) | (ps[4])) | ((ps[1]) | (ps[5]))) & (Areg[0])) & (Breg[1])) & (Preg[1])))) | ((((((ps[2]) | (ps[4])) | ((ps[1]) | (ps[5]))) & (Areg[0])) & (Breg[2])) & (Preg[2])))))));
    assign ready = ((~((_192_))));
    assign resultBus[0] = (Areg[0]);
    assign resultBus[1] = (Areg[1]);
    assign resultBus[2] = (Areg[2]);
    assign resultBus[3] = (Areg[3]);
    assign resultBus[4] = (Preg[0]);
    assign resultBus[5] = (Preg[1]);
    assign resultBus[6] = (Preg[2]);
    assign resultBus[7] = (Preg[3]);

endmodule