module Mult_Combinational_Sorted(
    input [3:0] ABus, BBus,
    input [3:0] Areg, Breg, Preg,
    input [5:1] ps,
    input _192_, start,

    output _193_, _024_, 
    output [3:0] _000_, _001_, _002_,
    output ready,
    output [7:0] resultBus
);

//   wire [3:0] _000_;
//   wire [3:0] _001_;
//   wire [3:0] _002_;
  wire _003_;
  wire _004_;
  wire _005_;
  wire _006_;
  wire _007_;
  wire _008_;
  wire _009_;
  wire _010_;
  wire _011_;
  wire _012_;
  wire _013_;
  wire _014_;
  wire _015_;
  wire _016_;
  wire _017_;
  wire _018_;
  wire _019_;
  wire _020_;
  wire _021_;
  wire _022_;
  wire _023_;
//   wire _024_;
  wire _025_;
  wire _026_;
  wire _027_;
  wire _028_;
  wire _029_;
  wire _030_;
  wire _031_;
  wire _032_;
  wire _033_;
  wire _034_;
  wire _035_;
  wire _036_;
  wire _037_;
  wire _038_;
  wire _039_;
  wire _040_;
  wire _041_;
  wire _042_;
  wire _043_;
  wire _044_;
  wire _045_;
  wire _046_;
  wire _047_;
  wire _048_;
  wire _049_;
  wire _050_;
  wire _051_;
  wire _052_;
  wire _053_;
  wire _054_;
  wire _055_;
  wire _056_;
  wire _057_;
  wire _058_;
  wire _059_;
  wire _060_;
  wire _061_;
  wire _062_;
  wire _063_;
  wire _064_;
  wire _065_;
  wire _066_;
  wire _067_;
  wire _068_;
  wire _069_;
  wire _070_;
  wire _071_;
  wire _072_;
  wire _073_;
  wire _074_;
  wire _075_;
  wire _076_;
  wire _077_;
  wire _078_;
  wire _079_;
  wire _080_;
  wire _081_;
  wire _082_;
  wire _083_;
  wire _084_;
  wire _085_;
  wire _086_;
  wire _087_;
  wire _088_;
  wire _089_;
  wire _090_;
  wire _091_;
  wire _092_;
  wire _093_;
  wire _094_;
  wire _095_;
  wire _096_;
  wire _097_;
  wire _098_;
  wire _099_;
  wire _100_;
  wire _101_;
  wire _102_;
  wire _103_;
  wire _104_;
  wire _105_;
  wire _106_;
  wire _107_;
  wire _108_;
  wire _109_;
  wire _110_;
  wire _111_;
  wire _112_;
  wire _113_;
  wire _114_;
  wire _115_;
  wire _116_;
  wire _117_;
  wire _118_;
  wire _119_;
  wire _120_;
  wire _121_;
  wire _122_;
  wire _123_;
  wire _124_;
  wire _125_;
  wire _126_;
  wire _127_;
  wire _128_;
  wire _129_;
  wire _130_;
  wire _131_;
  wire _132_;
  wire _133_;
  wire _134_;
  wire _135_;
  wire _136_;
  wire _137_;
  wire _138_;
  wire _139_;
  wire _140_;
  wire _141_;
  wire _142_;
  wire _143_;
  wire _144_;
  wire _145_;
  wire _146_;
  wire _147_;
  wire _148_;
  wire _149_;
  wire _150_;
  wire _151_;
  wire _152_;
  wire _153_;
  wire _154_;
  wire _155_;
  wire _156_;
  wire _157_;
  wire _158_;
  wire _159_;
  wire _160_;
  wire _161_;
  wire _162_;
  wire _163_;
  wire _164_;
  wire _165_;
  wire _166_;
  wire _167_;
  wire _168_;
  wire _169_;
  wire _170_;
  wire _171_;
  wire _172_;
  wire _173_;
  wire _174_;
  wire _175_;
  wire _176_;
  wire _177_;
  wire _178_;
  wire _179_;
  wire _180_;
  wire _181_;
  wire _182_;
  wire _183_;
  wire _184_;
  wire _185_;
  wire _186_;
  wire _187_;
  wire _188_;
  wire _189_;
  wire _190_;
  wire _191_;
  //wire _192_;
  //wire _193_;
  wire A0;
  //input [3:0] ABus;
  //wire [3:0] Areg;
  //input [3:0] BBus;
  //wire [3:0] Breg;
  //wire [3:0] Preg;
  //input clk;
  wire initP;
  wire loadA;
  wire loadB;
  //wire [5:0] ps;
  wire ps_0;
//   output ready;
//   output [7:0] resultBus;
  //input rst;
  //input start;

  assign A0 = Areg[0];
  assign initP = ps[3];
  assign loadA = ps[3];
  assign loadB = ps[3];
  assign resultBus = { Preg, Areg };
  assign _109_ = start;
  assign _129_ = Preg[0];
  assign _165_ = ps[4];
  assign _182_ = ps[5];
  assign _062_ = ps[1];
  assign _071_ = ps[2];
  assign _095_ = Breg[1];
  assign _101_ = Areg[0];
  assign _103_ = Preg[1];
  assign _104_ = Breg[0];
  assign _105_ = ps[3];
  assign _107_ = Preg[2];
  assign _108_ = Breg[2];
  assign _113_ = Breg[3];
  assign _114_ = Preg[3];
  assign _134_ = BBus[0];
  assign _138_ = BBus[1];
  assign _142_ = BBus[2];
  assign _146_ = BBus[3];
  assign _150_ = Areg[1];
  assign _153_ = ABus[0];
  assign _157_ = Areg[2];
  assign _160_ = ABus[1];
  assign _164_ = Areg[3];
  assign _167_ = ABus[2];
  assign _173_ = ABus[3];
  assign _179_ = _192_;

NOT _194_(_165_, _110_);
OR _195_(_179_, _109_, _112_);
AND _196_(_112_, _110_, _051_);
NOT _197_(_179_, _102_);
NOT _198_(_182_, _115_);
NOT _199_(_062_, _116_);
AND _200_(_116_, _115_, _117_);
NOT _201_(_071_, _118_);
AND _202_(_118_, _110_, _119_);
AND _203_(_119_, _117_, _120_);
OR _204_(_062_, _182_, _122_);
OR _205_(_071_, _165_, _123_);
OR _206_(_123_, _122_, _124_);
AND _207_(_124_, _101_, _125_);
AND _208_(_125_, _104_, _126_);
AND _209_(_126_, _129_, _127_);
NOT _210_(_127_, _128_);
NOT _211_(_103_, _130_);
NOT _212_(_095_, _131_);
NOT _213_(_101_, _133_);
OR _214_(_120_, _133_, _135_);
OR _215_(_135_, _131_, _137_);
AND _216_(_137_, _130_, _139_);
AND _217_(_125_, _095_, _141_);
AND _218_(_141_, _103_, _143_);
OR _219_(_143_, _139_, _145_);
OR _220_(_145_, _128_, _147_);
OR _221_(_141_, _103_, _149_);
OR _222_(_137_, _130_, _151_);
AND _223_(_151_, _149_, _152_);
OR _224_(_152_, _127_, _154_);
AND _225_(_154_, _147_, _156_);
OR _226_(_156_, _120_, _158_);
NOT _227_(_105_, _159_);
OR _228_(_124_, _129_, _161_);
AND _229_(_161_, _159_, _163_);
AND _230_(_163_, _158_, _106_);
AND _231_(_152_, _127_, _166_);
OR _232_(_166_, _143_, _168_);
AND _233_(_125_, _108_, _170_);
AND _234_(_170_, _107_, _171_);
NOT _235_(_171_, _172_);
OR _236_(_170_, _107_, _174_);
AND _237_(_174_, _172_, _176_);
OR _238_(_176_, _168_, _178_);
AND _239_(_147_, _151_, _180_);
NOT _240_(_176_, _181_);
OR _241_(_181_, _180_, _183_);
AND _242_(_183_, _178_, _184_);
OR _243_(_184_, _120_, _185_);
OR _244_(_124_, _103_, _186_);
AND _245_(_186_, _159_, _187_);
AND _246_(_187_, _185_, _111_);
AND _247_(_183_, _172_, _188_);
AND _248_(_125_, _113_, _189_);
OR _249_(_189_, _114_, _190_);
AND _250_(_189_, _114_, _191_);
NOT _251_(_191_, _052_);
AND _252_(_052_, _190_, _053_);
NOT _253_(_053_, _054_);
OR _254_(_054_, _188_, _055_);
AND _255_(_176_, _168_, _056_);
OR _256_(_056_, _171_, _057_);
OR _257_(_053_, _057_, _058_);
AND _258_(_058_, _055_, _059_);
OR _259_(_059_, _120_, _060_);
OR _260_(_124_, _107_, _061_);
AND _261_(_061_, _159_, _063_);
AND _262_(_063_, _060_, _121_);
AND _263_(_053_, _057_, _064_);
OR _264_(_191_, _120_, _065_);
OR _265_(_065_, _064_, _066_);
OR _266_(_124_, _114_, _067_);
AND _267_(_067_, _159_, _068_);
AND _268_(_068_, _066_, _132_);
OR _269_(_105_, _104_, _069_);
OR _270_(_134_, _159_, _070_);
AND _271_(_070_, _069_, _136_);
OR _272_(_105_, _095_, _072_);
OR _273_(_138_, _159_, _073_);
AND _274_(_073_, _072_, _140_);
OR _275_(_108_, _105_, _074_);
OR _276_(_142_, _159_, _075_);
AND _277_(_075_, _074_, _144_);
OR _278_(_113_, _105_, _076_);
OR _279_(_146_, _159_, _077_);
AND _280_(_077_, _076_, _148_);
AND _281_(_120_, _101_, _078_);
AND _282_(_124_, _150_, _079_);
OR _283_(_079_, _078_, _080_);
AND _284_(_080_, _159_, _081_);
AND _285_(_153_, _105_, _082_);
OR _286_(_082_, _081_, _155_);
AND _287_(_120_, _150_, _083_);
AND _288_(_124_, _157_, _084_);
OR _289_(_084_, _083_, _085_);
AND _290_(_085_, _159_, _086_);
AND _291_(_160_, _105_, _087_);
OR _292_(_087_, _086_, _162_);
AND _293_(_120_, _157_, _088_);
AND _294_(_124_, _164_, _089_);
OR _295_(_089_, _088_, _090_);
AND _296_(_090_, _159_, _091_);
AND _297_(_167_, _105_, _092_);
OR _298_(_092_, _091_, _169_);
OR _299_(_173_, _159_, _093_);
OR _300_(_126_, _129_, _094_);
AND _301_(_128_, _124_, _096_);
AND _302_(_096_, _094_, _097_);
AND _303_(_120_, _164_, _098_);
OR _304_(_098_, _105_, _099_);
OR _305_(_099_, _097_, _100_);
AND _306_(_100_, _093_, _175_);
AND _307_(_102_, _109_, _177_);


assign _193_ = _051_;
assign ready = ps_0;
assign ps_0 = _102_;
assign _002_[0] = _106_;
assign _002_[1] = _111_;
assign _002_[2] = _121_;
assign _002_[3] = _132_;
assign _001_[0] = _136_;
assign _001_[1] = _140_;
assign _001_[2] = _144_;
assign _001_[3] = _148_;
assign _000_[0] = _155_;
assign _000_[1] = _162_;
assign _000_[2] = _169_;
assign _000_[3] = _175_;
assign _024_ = _177_;

endmodule
